--fsm de melay, vhdl comportementale

library IEEE;
use IEEE.STD_LOGIC_1164.all;

entity mealy is
    port(clk    : in  STD_LOGIC;
         reset  : in  STD_LOGIC;
         input  : in  STD_LOGIC;
         output : out STD_LOGIC);
end;

architecture behavioral of mealy is
    type state_type is (s0, s1, s2, s3, s4, s5, s6);
    signal curr_state, next_state : state_type;
begin
    process(clk, reset)
    begin
        if (reset = '1') then
            curr_state <= s0;
        elsif (rising_edge(clk)) then
            curr_state <= next_state;
        end if;
    end process;

    process(curr_state, input)
    begin
        case curr_state is
            when s0 => -- a
                if (input = '0') then
                    output <= '0';
                    next_state <= s1;
                else
                    output <= '0';
                    next_state <= s2;
                end if;

            when s1 => -- b
				if (input = '0') then
                    output <= '0';
                    next_state <= s3;
                else
                    output <= '0';
                    next_state <= s4;
                end if;			
			
			when s2 => -- c
				if (input = '0') then
                    output <= '0';
                    next_state <= s5;
                else
                    output <= '0';
                    next_state <= s6;
                end if;
			
			when s3 => -- d	
				if (input = '0') then
                    output <= '0';
                    next_state <= s3;
                else
                    output <= '0';
                    next_state <= s4;
                end if;
			
			when s4 => -- e			
				if (input = '0') then
                    output <= '0';
                    next_state <= s5;
                else
                    output <= '1';
                    next_state <= s6;
                end if;
			
			when s5 => -- f			
				if (input = '0') then
                    output <= '0';
                    next_state <= s3;
                else
                    output <= '0';
                    next_state <= s4;
                end if;
			
			when s6 => -- g			
				if (input = '0') then
                    output <= '1';
                    next_state <= s5;
                else
                    output <= '0';
                    next_state <= s6;
                end if;
			
        end case;
    end process;
end;